//========================================================================
// DFFR_GL-test
//========================================================================

`include "ece2300/ece2300-test.v"

// ece2300-lint
`include "lab3/DFFR_GL.v"

module Top();

  //----------------------------------------------------------------------
  // Setup
  //----------------------------------------------------------------------

  CombinationalTestUtils t();

  //----------------------------------------------------------------------
  // Instantiate design under test
  //----------------------------------------------------------------------

  logic clk;
  logic rst;
  logic d;
  logic q;

  DFFR_GL dff
  (
    .clk (clk),
    .rst (rst),
    .d   (d),
    .q   (q)
  );

  //----------------------------------------------------------------------
  // Include test cases
  //----------------------------------------------------------------------

  `include "lab3/test/DFFR-test-cases.v"

endmodule

