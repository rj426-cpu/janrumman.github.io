//========================================================================
// BinaryToSevenSegUnopt_GL-test
//========================================================================

`include "ece2300/ece2300-test.v"

// ece2300-lint
`include "lab1/BinaryToSevenSegUnopt_GL.v"

module Top();

  //----------------------------------------------------------------------
  // Setup
  //----------------------------------------------------------------------

  CombinationalTestUtils t();

  //----------------------------------------------------------------------
  // Instantiate design under test
  //----------------------------------------------------------------------

  logic [3:0] in;
  logic [6:0] seg;

  BinaryToSevenSegUnopt_GL dut
  (
    .in  (in),
    .seg (seg)
  );

  //----------------------------------------------------------------------
  // Include test cases
  //----------------------------------------------------------------------

  `include "lab1/test/BinaryToSevenSeg-test-cases.v"

endmodule

