//========================================================================
// ImmGen_RTL-test
//========================================================================

`include "ece2300/ece2300-test.v"

// ece2300-lint
`include "lab4/ImmGen_RTL.v"

module Top();

  //----------------------------------------------------------------------
  // Setup
  //----------------------------------------------------------------------

  CombinationalTestUtils t();

  //----------------------------------------------------------------------
  // Instantiate design under test
  //----------------------------------------------------------------------

  logic [31:0] inst;
  logic  [1:0] imm_type;
  logic [31:0] imm;

  ImmGen_RTL dut
  (
    .inst     (inst),
    .imm_type (imm_type),
    .imm      (imm)
  );

  //----------------------------------------------------------------------
  // check
  //----------------------------------------------------------------------
  // We set the inputs, wait 8 tau, check the outputs, wait 2 tau. Each
  // check will take a total of 10 tau.

  task check
  (
    input logic [31:0] inst_,
    input logic  [1:0] imm_type_,
    input logic [31:0] imm_
  );
    if ( !t.failed ) begin
      t.num_checks += 1;

      inst     = inst_;
      imm_type = imm_type_;

      #8;

      if ( t.n != 0 )
        $display( "%3d: %h %d > %h", t.cycles, inst, imm_type, imm );

      `ECE2300_CHECK_EQ( imm, imm_ );

      #2;

    end
  endtask

  //----------------------------------------------------------------------
  // test_case_1_basic
  //----------------------------------------------------------------------

  task test_case_1_basic();
    t.test_case_begin( "test_case_1_basic" );

    //     inst           imm_type imm
    check( 32'h0000_0000, 0,       32'h0000_0000 );
    check( 32'h0000_0000, 1,       32'h0000_0000 );
    check( 32'h0000_0000, 2,       32'h0000_0000 );
    check( 32'h0000_0000, 3,       32'h0000_0000 );

    t.test_case_end();
  endtask

  //----------------------------------------------------------------------
  // test_case_2_directed_i_type
  //----------------------------------------------------------------------

  task test_case_2_directed_i_type();
    t.test_case_begin( "test_case_2_directed_i_type" );

    //         **** **** ****                                                           **** **** ****
    check( 32'b0000_0000_0000_0000_0000_0000_0000_0000, 0, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0001_0000_0000_0000_0000_0000, 0, 32'b0000_0000_0000_0000_0000_0000_0000_0001 );
    check( 32'b0101_0101_0101_0000_0000_0000_0000_0000, 0, 32'b0000_0000_0000_0000_0000_0101_0101_0101 );
    check( 32'b0110_1001_1111_0000_0000_0000_0000_0000, 0, 32'b0000_0000_0000_0000_0000_0110_1001_1111 );
    check( 32'b1000_0000_0000_0000_0000_0000_0000_0000, 0, 32'b1111_1111_1111_1111_1111_1000_0000_0000 );

    check( 32'b0000_0000_0000_1111_1111_1111_1111_1111, 0, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0001_1111_1111_1111_1111_1111, 0, 32'b0000_0000_0000_0000_0000_0000_0000_0001 );
    check( 32'b0101_0101_0101_1111_1111_1111_1111_1111, 0, 32'b0000_0000_0000_0000_0000_0101_0101_0101 );
    check( 32'b0110_1001_1111_1111_1111_1111_1111_1111, 0, 32'b0000_0000_0000_0000_0000_0110_1001_1111 );
    check( 32'b1000_0000_0000_1111_1111_1111_1111_1111, 0, 32'b1111_1111_1111_1111_1111_1000_0000_0000 );

    t.test_case_end();
  endtask

  //----------------------------------------------------------------------
  // test_case_3_directed_s_type
  //----------------------------------------------------------------------

  task test_case_3_directed_s_type();
    t.test_case_begin( "test_case_3_directed_s_type" );

    //         **** ***                 **** *                                          **** **** ****
    check( 32'b0000_0000_0000_0000_0000_0000_0000_0000, 1, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0000_0000_0000_0000_1000_0000, 1, 32'b0000_0000_0000_0000_0000_0000_0000_0001 );
    check( 32'b0010_1010_0000_0000_0000_1010_1000_0000, 1, 32'b0000_0000_0000_0000_0000_0010_1011_0101 );
    check( 32'b0110_1010_0000_0000_0000_1111_1000_0000, 1, 32'b0000_0000_0000_0000_0000_0110_1011_1111 );
    check( 32'b1000_0000_0000_0000_0000_0000_0000_0000, 1, 32'b1111_1111_1111_1111_1111_1000_0000_0000 );

    check( 32'b0000_0001_1111_1111_1111_0000_0111_1111, 1, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0001_1111_1111_1111_0000_1111_1111, 1, 32'b0000_0000_0000_0000_0000_0000_0000_0001 );
    check( 32'b0010_1011_1111_1111_1111_1010_1111_1111, 1, 32'b0000_0000_0000_0000_0000_0010_1011_0101 );
    check( 32'b0110_1011_1111_1111_1111_1111_1111_1111, 1, 32'b0000_0000_0000_0000_0000_0110_1011_1111 );
    check( 32'b1000_0001_1111_1111_1111_0000_0111_1111, 1, 32'b1111_1111_1111_1111_1111_1000_0000_0000 );

    t.test_case_end();
  endtask

  //----------------------------------------------------------------------
  // test_case_4_directed_j_type
  //----------------------------------------------------------------------

  task test_case_4_directed_j_type();
    t.test_case_begin( "test_case_4_directed_j_type" );

    //         abbb bbbb bbbc dddd dddd                                     a dddd dddd cbbb bbbb bbb0
    check( 32'b0000_0000_0000_0000_0000_0000_0000_0000, 2, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0010_0000_0000_0000_0000_0000, 2, 32'b0000_0000_0000_0000_0000_0000_0000_0010 );
    check( 32'b0010_1010_1011_1010_1010_0000_0000_0000, 2, 32'b0000_0000_0000_1010_1010_1010_1010_1010 );
    check( 32'b1000_0000_0000_0000_0000_0000_0000_0000, 2, 32'b1111_1111_1111_0000_0000_0000_0000_0000 );

    check( 32'b0000_0000_0000_0000_0000_1111_1111_1111, 2, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0010_0000_0000_1111_1111_1111, 2, 32'b0000_0000_0000_0000_0000_0000_0000_0010 );
    check( 32'b0010_1010_1011_1010_1010_1111_1111_1111, 2, 32'b0000_0000_0000_1010_1010_1010_1010_1010 );
    check( 32'b1000_0000_0000_0000_0000_1111_1111_1111, 2, 32'b1111_1111_1111_0000_0000_0000_0000_0000 );

    t.test_case_end();
  endtask

  //----------------------------------------------------------------------
  // test_case_5_directed_b_type
  //----------------------------------------------------------------------

  task test_case_5_directed_b_type();
    t.test_case_begin( "test_case_5_directed_b_type" );

    //         abbb bbb                 dddd c                                        a cbbb bbbd ddd0
    check( 32'b0000_0000_0000_0000_0000_0000_0000_0000, 3, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0000_0000_0000_0001_0000_0000, 3, 32'b0000_0000_0000_0000_0000_0000_0000_0010 );
    check( 32'b0010_1010_0000_0000_0000_0101_1000_0000, 3, 32'b0000_0000_0000_0000_0000_1010_1010_1010 );
    check( 32'b1000_0000_0000_0000_0000_0000_0000_0000, 3, 32'b1111_1111_1111_1111_1111_0000_0000_0000 );

    check( 32'b0000_0001_1111_1111_1111_0000_0111_1111, 3, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0001_1111_1111_1111_0001_0111_1111, 3, 32'b0000_0000_0000_0000_0000_0000_0000_0010 );
    check( 32'b0010_1011_1111_1111_1111_0101_1111_1111, 3, 32'b0000_0000_0000_0000_0000_1010_1010_1010 );
    check( 32'b1000_0001_1111_1111_1111_0000_0111_1111, 3, 32'b1111_1111_1111_1111_1111_0000_0000_0000 );

    t.test_case_end();
  endtask

  //----------------------------------------------------------------------
  // test_case_6_xprop
  //----------------------------------------------------------------------

  task test_case_6_xprop();
    t.test_case_begin( "test_case_6_xprop" );

    //     inst imm_type imm
    check( 'x,  'x,      'x );

    t.test_case_end();
  endtask

  //----------------------------------------------------------------------
  // main
  //----------------------------------------------------------------------

  initial begin
    t.test_bench_begin();

    if ((t.n <= 0) || (t.n == 1)) test_case_1_basic();
    if ((t.n <= 0) || (t.n == 2)) test_case_2_directed_i_type();
    if ((t.n <= 0) || (t.n == 3)) test_case_3_directed_s_type();
    if ((t.n <= 0) || (t.n == 4)) test_case_4_directed_j_type();
    if ((t.n <= 0) || (t.n == 5)) test_case_5_directed_b_type();
    if ((t.n <= 0) || (t.n == 6)) test_case_6_xprop();

    t.test_bench_end();
  end

endmodule

