//========================================================================
// Multiplier_2x8b_GL-test
//========================================================================

`include "ece2300/ece2300-test.v"

// ece2300-lint
`include "lab2/Multiplier_2x16b_GL.v"

module Top();

  //----------------------------------------------------------------------
  // Setup
  //----------------------------------------------------------------------

  CombinationalTestUtils t();

  //----------------------------------------------------------------------
  // Instantiate design under test
  //----------------------------------------------------------------------

  logic [15:0] in0;
  logic  [1:0] in1;
  logic [15:0] prod;

  Multiplier_2x16b_GL dut
  (
    .in0  (in0),
    .in1  (in1),
    .prod (prod)
  );

  //----------------------------------------------------------------------
  // Include test cases
  //----------------------------------------------------------------------

  `include "lab2/test/Multiplier_2x16b-test-cases.v"

endmodule

