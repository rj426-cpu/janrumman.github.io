//========================================================================
// DisplayOpt_GL-test
//========================================================================

`include "ece2300/ece2300-test.v"

// ece2300-lint
`include "lab1/DisplayOpt_GL.v"

module Top();

  //----------------------------------------------------------------------
  // Setup
  //----------------------------------------------------------------------

  CombinationalTestUtils t();

  //----------------------------------------------------------------------
  // Instantiate design under test
  //----------------------------------------------------------------------

  logic [4:0] in;
  logic [6:0] seg_tens;
  logic [6:0] seg_ones;

  DisplayOpt_GL dut
  (
    .in       (in),
    .seg_tens (seg_tens),
    .seg_ones (seg_ones)
  );

  //----------------------------------------------------------------------
  // Include test cases
  //----------------------------------------------------------------------

  `include "lab1/test/Display-test-cases.v"

endmodule

