//========================================================================
// Register_16b_RTL-test
//========================================================================

`include "ece2300/ece2300-test.v"

// ece2300-lint
`include "lab3/Register_16b_RTL.v"

module Top();

  //----------------------------------------------------------------------
  // Setup
  //----------------------------------------------------------------------

  logic clk;
  logic rst_foo;

  TestUtilsClkRst t
  (
    .clk (clk),
    .rst (rst_foo)
  );

  //----------------------------------------------------------------------
  // Instantiate design under test
  //----------------------------------------------------------------------

  logic        rst;
  logic        en;
  logic [15:0] d;
  logic [15:0] q;

  Register_16b_RTL register
  (
    .clk (clk),
    .rst (rst | rst_foo),
    .en  (en),
    .d   (d),
    .q   (q)
  );

  //----------------------------------------------------------------------
  // Include test cases
  //----------------------------------------------------------------------

  `include "lab3/test/Register_16b-test-cases.v"

endmodule

