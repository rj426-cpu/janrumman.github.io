//========================================================================
// AdderCarrySelect_16b_GL-test
//========================================================================

`include "ece2300/ece2300-test.v"

// ece2300-lint
`include "lab2/AdderCarrySelect_16b_GL.v"

module Top();

  //----------------------------------------------------------------------
  // Setup
  //----------------------------------------------------------------------

  CombinationalTestUtils t();

  //----------------------------------------------------------------------
  // Instantiate design under test
  //----------------------------------------------------------------------

  logic [15:0] in0;
  logic [15:0] in1;
  logic        cin;
  logic        cout;
  logic [15:0] sum;

  AdderCarrySelect_16b_GL dut
  (
    .in0  (in0),
    .in1  (in1),
    .cin  (cin),
    .cout (cout),
    .sum  (sum)
  );

  //----------------------------------------------------------------------
  // Include test cases
  //----------------------------------------------------------------------

  `include "lab2/test/Adder_16b-test-cases.v"

endmodule

